class sequencer extends component_base;
	function new (string name, component_base parent);
	    this.name = name;
	    this.parent = parent;
	  endfunction
endclass
